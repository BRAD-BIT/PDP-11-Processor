LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY my_adder IS
    PORT( a,b,cin : IN  std_logic; s,cout : OUT  std_logic);
END ENTITY my_adder;

ARCHITECTURE behav OF my_adder IS
BEGIN
        PROCESS (a,b,cin)     
	BEGIN
        s <= a XOR b XOR cin;
        cout <= (a AND b) or (cin AND (a XOR b));
	END PROCESS;
END behav;
